package ahb_master_pkg;
	import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "ahb_trans.sv"
    `include "ahb_sequence.sv"
    `include "ahb_driver.sv"
    `include "ahb_sqr.sv"
    `include "ahb_monitor.sv"
    `include "ahb_agt.sv"
    
endpackage