package apb_slave_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "apb_trans.sv"
	`include "apb_sequence.sv"
	`include "apb_driver.sv"
	`include "apb_sqr.sv"
	`include "apb_monitor.sv"
	`include "apb_agt.sv"
	
endpackage